module helloworld();
	initial begin 
		$display ("My name is Janani P Srinivasan and I start the course today 05/04/2025!");
	end

endmodule
