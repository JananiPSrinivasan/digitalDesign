`timescale 1ns/1ns

module nbitdecoder_tb();
endmodule