module (
    input clk,
    input rst,
    input reg [3:0] d,
    output q
);
    
endmodule